module LEGz_Architecture (clk, rst, Output_1, Output_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [7:0] Output_1;
  output  wire [7:0] Output_2;

  TC_Counter # (.UUID(64'd2124775489427933008 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_0 (.clk(clk), .rst(rst), .save(wire_56), .in(wire_13), .out(wire_32));
  TC_Splitter8 # (.UUID(64'd4551787757548942711 ^ UUID)) Splitter8_1 (.in({{7{1'b0}}, wire_30 }), .out0(wire_74), .out1(wire_27), .out2(wire_71), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3796524371277023761 ^ UUID)) Decoder3_2 (.dis(wire_2), .sel0(wire_74), .sel1(wire_27), .sel2(wire_71), .out0(wire_81), .out1(wire_62), .out2(wire_64), .out3(wire_18), .out4(wire_65), .out5(wire_59), .out6(wire_7), .out7(wire_85));
  TC_Switch # (.UUID(64'd2063467048664777668 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_52), .in(wire_37), .out(wire_14_7));
  TC_Switch # (.UUID(64'd3378363622096012442 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_3), .in(wire_24), .out(wire_14_6));
  TC_Switch # (.UUID(64'd4371098375043748744 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_16), .in(wire_11), .out(wire_14_5));
  TC_Switch # (.UUID(64'd238512083288038597 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_25), .in(wire_29), .out(wire_14_4));
  TC_Switch # (.UUID(64'd64626453180078677 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_44), .in(wire_57), .out(wire_14_3));
  TC_Switch # (.UUID(64'd317325102133445192 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_87), .in(wire_31), .out(wire_14_2));
  TC_Switch # (.UUID(64'd214230785942808532 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_83), .in(wire_32), .out(wire_14_0));
  TC_Switch # (.UUID(64'd2210798626195217718 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_50), .in({{7{1'b0}}, wire_55 }), .out(wire_14_1));
  TC_Switch # (.UUID(64'd433540470023572044 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_70), .in(wire_24), .out(wire_23_2));
  TC_Switch # (.UUID(64'd2763545113978640643 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_17), .in(wire_11), .out(wire_23_3));
  TC_Switch # (.UUID(64'd2074149251288325490 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_20), .in(wire_29), .out(wire_23_4));
  TC_Switch # (.UUID(64'd2425319554433863854 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_6), .in(wire_57), .out(wire_23_5));
  TC_Switch # (.UUID(64'd2696410939672307921 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_61), .in(wire_31), .out(wire_23_6));
  TC_Switch # (.UUID(64'd3912814052070262056 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_67), .in(wire_32), .out(wire_23_7));
  TC_Switch # (.UUID(64'd3559162101923647238 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_46), .in({{7{1'b0}}, wire_55 }), .out(wire_23_8));
  TC_Splitter8 # (.UUID(64'd532206217823046164 ^ UUID)) Splitter8_18 (.in({{7{1'b0}}, wire_5 }), .out0(wire_26), .out1(wire_79), .out2(wire_76), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd1155637373704071995 ^ UUID)) Decoder3_19 (.dis(wire_38), .sel0(wire_26), .sel1(wire_79), .sel2(wire_76), .out0(wire_21), .out1(wire_70), .out2(wire_17), .out3(wire_20), .out4(wire_6), .out5(wire_61), .out6(wire_67), .out7(wire_46));
  TC_Splitter8 # (.UUID(64'd2397136406627350888 ^ UUID)) Splitter8_20 (.in({{7{1'b0}}, wire_4 }), .out0(wire_73), .out1(wire_34), .out2(wire_42), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2812330477263231948 ^ UUID)) Decoder3_21 (.dis(wire_15), .sel0(wire_73), .sel1(wire_34), .sel2(wire_42), .out0(wire_52), .out1(wire_3), .out2(wire_16), .out3(wire_25), .out4(wire_44), .out5(wire_87), .out6(wire_83), .out7(wire_50));
  TC_Switch # (.UUID(64'd2727240096060367728 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_22 (.en(wire_25), .in(wire_25), .out(wire_40_0));
  TC_Switch # (.UUID(64'd2049181701106783432 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_23 (.en(wire_44), .in(wire_44), .out(wire_9_0));
  TC_Switch # (.UUID(64'd2482488626744003376 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_24 (.en(wire_87), .in(wire_87), .out(wire_88_0));
  TC_Switch # (.UUID(64'd1958765381208861188 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_25 (.en(wire_20), .in(wire_20), .out(wire_40_1));
  TC_Switch # (.UUID(64'd3924109062529388782 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_26 (.en(wire_6), .in(wire_6), .out(wire_9_1));
  TC_Switch # (.UUID(64'd632104071497708010 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_27 (.en(wire_61), .in(wire_61), .out(wire_88_1));
  TC_Switch # (.UUID(64'd3061836083092996367 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_7), .in(wire_48), .out(wire_13_0));
  TC_Switch # (.UUID(64'd618709936422461351 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_15), .in({{7{1'b0}}, wire_4 }), .out(wire_14_8));
  TC_Switch # (.UUID(64'd1628120986469259568 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_38), .in({{7{1'b0}}, wire_5 }), .out(wire_23_0));
  TC_Switch # (.UUID(64'd3004464700760938994 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_10), .in({{7{1'b0}}, wire_30 }), .out(wire_84));
  TC_Switch # (.UUID(64'd2943121197558932545 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_32 (.en(wire_7), .in(wire_7), .out(wire_56_0));
  TC_Switch # (.UUID(64'd2529615440270560801 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_21), .in(wire_37), .out(wire_23_1));
  TC_Switch # (.UUID(64'd3239767307943638156 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_66), .in(wire_66), .out(wire_10_2));
  TC_Ram # (.UUID(64'd2888211812749069423 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_35 (.clk(clk), .rst(rst), .load(wire_49), .save(wire_1), .address({{24{1'b0}}, wire_78 }), .in0({{56{1'b0}}, wire_23 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_68), .out1(), .out2(), .out3());
  TC_Register # (.UUID(64'd4589497095347758610 ^ UUID), .BIT_WIDTH(64'd8)) Register8_36 (.clk(clk), .rst(rst), .load(wire_47), .save(wire_81), .in(wire_48), .out(wire_37));
  TC_Register # (.UUID(64'd4196636957227629122 ^ UUID), .BIT_WIDTH(64'd8)) Register8_37 (.clk(clk), .rst(rst), .load(wire_43), .save(wire_62), .in(wire_48), .out(wire_24));
  TC_Register # (.UUID(64'd2337026380131603269 ^ UUID), .BIT_WIDTH(64'd8)) Register8_38 (.clk(clk), .rst(rst), .load(wire_72), .save(wire_64), .in(wire_48), .out(wire_11));
  TC_Register # (.UUID(64'd4391459169503373385 ^ UUID), .BIT_WIDTH(64'd8)) Register8_39 (.clk(clk), .rst(rst), .load(wire_9), .save(wire_65), .in(wire_48), .out(wire_57));
  TC_Register # (.UUID(64'd542874102567414615 ^ UUID), .BIT_WIDTH(64'd8)) Register8_40 (.clk(clk), .rst(rst), .load(wire_88), .save(wire_59), .in(wire_48), .out(wire_31));
  TC_Switch # (.UUID(64'd4032239855974584733 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_41 (.en(wire_1), .in(wire_60), .out(wire_78_0));
  TC_Switch # (.UUID(64'd4569436211148002821 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_42 (.en(wire_49), .in(wire_60), .out(wire_78_1));
  TC_Switch # (.UUID(64'd651672442968330745 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_43 (.en(wire_49), .in(wire_68[7:0]), .out(wire_22_0));
  TC_Switch # (.UUID(64'd1957120000915480017 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_12), .in(wire_14), .out(wire_39_0));
  TC_Mux # (.UUID(64'd503367712643433779 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_45 (.sel(wire_36), .in0(wire_84), .in1(wire_22), .out(wire_13_1));
  TC_Switch # (.UUID(64'd285289608810659520 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_46 (.en(wire_52), .in(wire_52), .out(wire_47_0));
  TC_Switch # (.UUID(64'd1149378019528028669 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_47 (.en(wire_21), .in(wire_21), .out(wire_47_1));
  TC_Switch # (.UUID(64'd4605667724210175680 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_48 (.en(wire_70), .in(wire_70), .out(wire_43_0));
  TC_Switch # (.UUID(64'd3394422510326288105 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_49 (.en(wire_3), .in(wire_3), .out(wire_43_1));
  TC_Switch # (.UUID(64'd4567104258324075038 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_50 (.en(wire_17), .in(wire_17), .out(wire_72_1));
  TC_Switch # (.UUID(64'd401433735891713226 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_51 (.en(wire_16), .in(wire_16), .out(wire_72_0));
  TC_Switch # (.UUID(64'd1483338896357059824 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_45), .in(wire_75), .out(wire_48_2));
  TC_Register # (.UUID(64'd1457531445102985096 ^ UUID), .BIT_WIDTH(64'd8)) Register8_53 (.clk(clk), .rst(rst), .load(wire_40), .save(wire_18), .in(wire_48), .out(wire_29));
  TC_Switch # (.UUID(64'd544989980592214467 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_63), .in(wire_19), .out(wire_39_1));
  TC_Switch # (.UUID(64'd3421564125831961817 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_55 (.en(wire_54), .in(wire_39), .out(wire_60_0));
  TC_Switch # (.UUID(64'd2237576448329743067 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_56 (.en(wire_77), .in(wire_33), .out(wire_48_3));
  TC_Switch # (.UUID(64'd4055037871993213722 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_57 (.en(wire_41), .in(wire_22), .out(wire_48_0));
  TC_Switch # (.UUID(64'd3415539481769456348 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_58 (.en(wire_80), .in(wire_80), .out(wire_10_0));
  TC_Switch # (.UUID(64'd101413649404046443 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_59 (.en(wire_86), .in(wire_48), .out(Output_2));
  TC_Switch # (.UUID(64'd2192670883954912709 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_60 (.en(wire_58), .in({{7{1'b0}}, wire_55 }), .out(Output_1));
  Comparatorz_zmz_Unsigned # (.UUID(64'd3039673388688779802 ^ UUID)) Comparatorz_zmz_Unsigned_61 (.clk(clk), .rst(rst), .Opcode({{7{1'b0}}, wire_28 }), .Input_1(wire_14), .Input_2(wire_23), .Output(wire_66));
  Stack # (.UUID(64'd3850316400058731886 ^ UUID)) Stack_62 (.clk(clk), .rst(rst), .POP(wire_69), .PUSH(wire_51), .VALUE(wire_60), .OUTPUT(wire_22_1));
  Storagez_Controller # (.UUID(64'd790116534102722917 ^ UUID)) Storagez_Controller_63 (.clk(clk), .rst(rst), .ControlBus({{7{1'b0}}, wire_28 }), .CurrentCounter(wire_32), .ReturnCounter(wire_60_1), .DisableDataBus(wire_35), .EnableRamAddress(wire_54), .Overwrite(wire_10_1), .STORE(wire_1), .LOAD(wire_49), .PUSH(wire_8), .MuxStorageOut(wire_82), .RemainderToStack(wire_63), .POP(wire_69), .EnableStorageOut(wire_53));
  LSL # (.UUID(64'd1376843152744323112 ^ UUID)) LSL_64 (.clk(clk), .rst(rst), .value(wire_23), .num_shift_4bit(wire_14), .\output (wire_75));
  Addressz_Busz_Controller # (.UUID(64'd310120577754861117 ^ UUID)) Addressz_Busz_Controller_65 (.clk(clk), .rst(rst), .OP_Code({{7{1'b0}}, wire_28 }), .IMMA(wire_15_1), .IMMB(wire_38_1), .IMMALL(wire_0), .LSL(wire_45), .LSR(wire_77));
  _1bz_buffersz_x4 # (.UUID(64'd86212022713044376 ^ UUID)) _1bz_buffersz_x4_66 (.clk(clk), .rst(rst), .Input1(wire_46), .Input2(1'd0), .Input3(1'd0), .Input4(wire_50), .Output1(wire_58_2), .Output2(wire_58_0), .Output3(wire_58_1), .Output4(wire_58_3));
  ALUz_zmz_LEG # (.UUID(64'd3446037741910496325 ^ UUID)) ALUz_zmz_LEG_67 (.clk(clk), .rst(rst), .Opcode({{7{1'b0}}, wire_28 }), .Input_1(wire_14), .Input_2(wire_23), .Output(wire_48_1), .Carry(wire_19));
  _1bz_buffersz_x4 # (.UUID(64'd2043273707421821908 ^ UUID)) _1bz_buffersz_x4_68 (.clk(clk), .rst(rst), .Input1(wire_8), .Input2(wire_53), .Input3(wire_82), .Input4(wire_63), .Output1(wire_51_0), .Output2(wire_41), .Output3(wire_36), .Output4(wire_51_1));
  _1bz_buffersz_x4 # (.UUID(64'd2914315711682501393 ^ UUID)) _1bz_buffersz_x4_69 (.clk(clk), .rst(rst), .Input1(wire_1), .Input2(wire_1), .Input3(wire_49), .Input4(wire_8), .Output1(wire_2_3), .Output2(wire_12_2), .Output3(wire_12_0), .Output4(wire_12_1));
  LSR # (.UUID(64'd505032913097474618 ^ UUID)) LSR_70 (.clk(clk), .rst(rst), .Value(wire_23), .\4bit_shift_num (wire_14), .OUT(wire_33));
  _1bz_buffersz_x2 # (.UUID(64'd3015520887090458698 ^ UUID)) _1bz_buffersz_x2_71 (.clk(clk), .rst(rst), .Input1(wire_10), .Input2(wire_10), .Output1(wire_56_1), .Output2(wire_2_0));
  _1bz_buffersz_x2 # (.UUID(64'd544146479927488242 ^ UUID)) _1bz_buffersz_x2_72 (.clk(clk), .rst(rst), .Input1(wire_0), .Input2(wire_0), .Output1(wire_15_0), .Output2(wire_38_0));
  _1bz_buffersz_x2 # (.UUID(64'd2995839097132858056 ^ UUID)) _1bz_buffersz_x2_73 (.clk(clk), .rst(rst), .Input1(wire_85), .Input2(1'd0), .Output1(wire_86), .Output2());
  _1bz_buffersz_x2 # (.UUID(64'd2738157904611306808 ^ UUID)) _1bz_buffersz_x2_74 (.clk(clk), .rst(rst), .Input1(wire_35), .Input2(wire_8), .Output1(wire_2_1), .Output2(wire_2_2));
  Comparatorz_zmz_Signed # (.UUID(64'd3192642732172097703 ^ UUID)) Comparatorz_zmz_Signed_75 (.clk(clk), .rst(rst), .Opcode({{7{1'b0}}, wire_28 }), .Input_1(wire_14), .Input_2(wire_23), .Output(wire_80));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_2_0;
  wire [0:0] wire_2_1;
  wire [0:0] wire_2_2;
  wire [0:0] wire_2_3;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  assign wire_4 = 0;
  wire [0:0] wire_5;
  assign wire_5 = 0;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_9_0;
  wire [0:0] wire_9_1;
  assign wire_9 = wire_9_0|wire_9_1;
  wire [0:0] wire_10;
  wire [0:0] wire_10_0;
  wire [0:0] wire_10_1;
  wire [0:0] wire_10_2;
  assign wire_10 = wire_10_0|wire_10_1|wire_10_2;
  wire [7:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_12_0;
  wire [0:0] wire_12_1;
  wire [0:0] wire_12_2;
  assign wire_12 = wire_12_0|wire_12_1|wire_12_2;
  wire [7:0] wire_13;
  wire [7:0] wire_13_0;
  wire [7:0] wire_13_1;
  assign wire_13 = wire_13_0|wire_13_1;
  wire [7:0] wire_14;
  wire [7:0] wire_14_0;
  wire [7:0] wire_14_1;
  wire [7:0] wire_14_2;
  wire [7:0] wire_14_3;
  wire [7:0] wire_14_4;
  wire [7:0] wire_14_5;
  wire [7:0] wire_14_6;
  wire [7:0] wire_14_7;
  wire [7:0] wire_14_8;
  assign wire_14 = wire_14_0|wire_14_1|wire_14_2|wire_14_3|wire_14_4|wire_14_5|wire_14_6|wire_14_7|wire_14_8;
  wire [0:0] wire_15;
  wire [0:0] wire_15_0;
  wire [0:0] wire_15_1;
  assign wire_15 = wire_15_0|wire_15_1;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [7:0] wire_22_0;
  wire [7:0] wire_22_1;
  assign wire_22 = wire_22_0|wire_22_1;
  wire [7:0] wire_23;
  wire [7:0] wire_23_0;
  wire [7:0] wire_23_1;
  wire [7:0] wire_23_2;
  wire [7:0] wire_23_3;
  wire [7:0] wire_23_4;
  wire [7:0] wire_23_5;
  wire [7:0] wire_23_6;
  wire [7:0] wire_23_7;
  wire [7:0] wire_23_8;
  assign wire_23 = wire_23_0|wire_23_1|wire_23_2|wire_23_3|wire_23_4|wire_23_5|wire_23_6|wire_23_7|wire_23_8;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  assign wire_28 = 0;
  wire [7:0] wire_29;
  wire [0:0] wire_30;
  assign wire_30 = 0;
  wire [7:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_38_0;
  wire [0:0] wire_38_1;
  assign wire_38 = wire_38_0|wire_38_1;
  wire [7:0] wire_39;
  wire [7:0] wire_39_0;
  wire [7:0] wire_39_1;
  assign wire_39 = wire_39_0|wire_39_1;
  wire [0:0] wire_40;
  wire [0:0] wire_40_0;
  wire [0:0] wire_40_1;
  assign wire_40 = wire_40_0|wire_40_1;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_43_0;
  wire [0:0] wire_43_1;
  assign wire_43 = wire_43_0|wire_43_1;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_47_0;
  wire [0:0] wire_47_1;
  assign wire_47 = wire_47_0|wire_47_1;
  wire [7:0] wire_48;
  wire [7:0] wire_48_0;
  wire [7:0] wire_48_1;
  wire [7:0] wire_48_2;
  wire [7:0] wire_48_3;
  assign wire_48 = wire_48_0|wire_48_1|wire_48_2|wire_48_3;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_51_0;
  wire [0:0] wire_51_1;
  assign wire_51 = wire_51_0|wire_51_1;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  assign wire_55 = 0;
  wire [0:0] wire_56;
  wire [0:0] wire_56_0;
  wire [0:0] wire_56_1;
  assign wire_56 = wire_56_0|wire_56_1;
  wire [7:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_58_0;
  wire [0:0] wire_58_1;
  wire [0:0] wire_58_2;
  wire [0:0] wire_58_3;
  assign wire_58 = wire_58_0|wire_58_1|wire_58_2|wire_58_3;
  wire [0:0] wire_59;
  wire [7:0] wire_60;
  wire [7:0] wire_60_0;
  wire [7:0] wire_60_1;
  assign wire_60 = wire_60_0|wire_60_1;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [63:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_72_0;
  wire [0:0] wire_72_1;
  assign wire_72 = wire_72_0|wire_72_1;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [7:0] wire_78;
  wire [7:0] wire_78_0;
  wire [7:0] wire_78_1;
  assign wire_78 = wire_78_0|wire_78_1;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_88_0;
  wire [0:0] wire_88_1;
  assign wire_88 = wire_88_0|wire_88_1;

endmodule
