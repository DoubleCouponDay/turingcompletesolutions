module Stack (clk, rst, POP, PUSH, VALUE, OUTPUT);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] POP;
  input  wire [0:0] PUSH;
  input  wire [7:0] VALUE;
  output  wire [7:0] OUTPUT;

  TC_Switch # (.UUID(64'd8301479748015613097 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_0 (.en(wire_5), .in(wire_12), .out(OUTPUT));
  TC_Register # (.UUID(64'd3792999861150587255 ^ UUID), .BIT_WIDTH(64'd8)) Register8_1 (.clk(clk), .rst(rst), .load(wire_8), .save(wire_49), .in(wire_3), .out(wire_12_14));
  TC_Register # (.UUID(64'd1058998454388883399 ^ UUID), .BIT_WIDTH(64'd8)) Register8_2 (.clk(clk), .rst(rst), .load(wire_41), .save(wire_51), .in(wire_3), .out(wire_12_13));
  TC_Register # (.UUID(64'd3634169620936557151 ^ UUID), .BIT_WIDTH(64'd8)) Register8_3 (.clk(clk), .rst(rst), .load(wire_59), .save(wire_37), .in(wire_3), .out(wire_12_12));
  TC_Register # (.UUID(64'd3787560344221118625 ^ UUID), .BIT_WIDTH(64'd8)) Register8_4 (.clk(clk), .rst(rst), .load(wire_53), .save(wire_21), .in(wire_3), .out(wire_12_11));
  TC_Register # (.UUID(64'd2413072079755975483 ^ UUID), .BIT_WIDTH(64'd8)) Register8_5 (.clk(clk), .rst(rst), .load(wire_23), .save(wire_42), .in(wire_3), .out(wire_12_10));
  TC_Register # (.UUID(64'd2548569033097971443 ^ UUID), .BIT_WIDTH(64'd8)) Register8_6 (.clk(clk), .rst(rst), .load(wire_56), .save(wire_48), .in(wire_3), .out(wire_12_9));
  TC_Register # (.UUID(64'd3394111936823370531 ^ UUID), .BIT_WIDTH(64'd8)) Register8_7 (.clk(clk), .rst(rst), .load(wire_57), .save(wire_18), .in(wire_3), .out(wire_12_4));
  TC_Splitter8 # (.UUID(64'd3792967820205480956 ^ UUID)) Splitter8_8 (.in(wire_33), .out0(wire_55), .out1(wire_61), .out2(wire_11), .out3(wire_34), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3681355771047358362 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_9 (.en(wire_7), .in(wire_32), .out(wire_49));
  TC_Switch # (.UUID(64'd2629695715771492218 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_10 (.en(wire_7), .in(wire_30), .out(wire_51));
  TC_Switch # (.UUID(64'd2486263146412058506 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(wire_10), .in(wire_1), .out(wire_59));
  TC_Switch # (.UUID(64'd1075832990892126228 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_12 (.en(wire_7), .in(wire_17), .out(wire_21));
  TC_Switch # (.UUID(64'd2576687253761336672 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_13 (.en(wire_7), .in(wire_40), .out(wire_42));
  TC_Switch # (.UUID(64'd1569695276672358489 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_7), .in(wire_4), .out(wire_48));
  TC_Switch # (.UUID(64'd1081270592699420271 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_15 (.en(wire_7), .in(wire_13), .out(wire_18));
  TC_Switch # (.UUID(64'd2107057030057130682 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_16 (.en(wire_10), .in(wire_17), .out(wire_53));
  TC_Switch # (.UUID(64'd4530925573592076500 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_10), .in(wire_40), .out(wire_23));
  TC_Switch # (.UUID(64'd3419148342944904523 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_18 (.en(wire_10), .in(wire_4), .out(wire_56));
  TC_Switch # (.UUID(64'd2586762651624420451 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_19 (.en(wire_10), .in(wire_13), .out(wire_57));
  TC_Switch # (.UUID(64'd851354254291366217 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_20 (.en(wire_10), .in(wire_32), .out(wire_8));
  TC_Switch # (.UUID(64'd1497549122964121087 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_21 (.en(wire_10), .in(wire_30), .out(wire_41));
  TC_Switch # (.UUID(64'd430849778933204556 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_22 (.en(wire_7), .in(wire_1), .out(wire_37));
  TC_Switch # (.UUID(64'd3795977666512523172 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_23 (.en(wire_5), .in(wire_5), .out(wire_10));
  TC_Switch # (.UUID(64'd4009430940610121027 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_24 (.en(wire_2), .in(wire_2), .out(wire_7));
  TC_Constant # (.UUID(64'd1489445187687683920 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hFF)) Constant8_25 (.out(wire_50));
  TC_Constant # (.UUID(64'd197535579952262412 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_26 (.out(wire_19));
  TC_Add # (.UUID(64'd1472804865791430980 ^ UUID), .BIT_WIDTH(64'd8)) Add8_27 (.in0(wire_9), .in1(wire_16), .ci(1'd0), .out(wire_14), .co());
  TC_Register # (.UUID(64'd963982926232964878 ^ UUID), .BIT_WIDTH(64'd8)) Register8_28 (.clk(clk), .rst(rst), .load(wire_22), .save(wire_22), .in(wire_14), .out(wire_9));
  TC_Switch # (.UUID(64'd3587542012384850459 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_5), .in(wire_50), .out(wire_16_0));
  TC_Switch # (.UUID(64'd4190922332537850963 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_2), .in(wire_19), .out(wire_16_1));
  TC_Switch # (.UUID(64'd1242448487826305409 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_31 (.en(wire_5), .in(wire_5), .out(wire_22_0));
  TC_Switch # (.UUID(64'd4015284971698115546 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_32 (.en(wire_2), .in(wire_2), .out(wire_22_1));
  TC_Mux # (.UUID(64'd1774473313025810126 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_33 (.sel(wire_2), .in0(wire_9), .in1(wire_14), .out(wire_33));
  TC_Register # (.UUID(64'd4538217995780326528 ^ UUID), .BIT_WIDTH(64'd8)) Register8_34 (.clk(clk), .rst(rst), .load(wire_25), .save(wire_43), .in(wire_3), .out(wire_12_6));
  TC_Register # (.UUID(64'd427235039069631583 ^ UUID), .BIT_WIDTH(64'd8)) Register8_35 (.clk(clk), .rst(rst), .load(wire_46), .save(wire_60), .in(wire_3), .out(wire_12_8));
  TC_Register # (.UUID(64'd1332592916367643629 ^ UUID), .BIT_WIDTH(64'd8)) Register8_36 (.clk(clk), .rst(rst), .load(wire_58), .save(wire_54), .in(wire_3), .out(wire_12_3));
  TC_Register # (.UUID(64'd4057818994473822135 ^ UUID), .BIT_WIDTH(64'd8)) Register8_37 (.clk(clk), .rst(rst), .load(wire_39), .save(wire_38), .in(wire_3), .out(wire_12_1));
  TC_Switch # (.UUID(64'd725527960586846217 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_38 (.en(wire_10), .in(wire_24), .out(wire_25));
  TC_Switch # (.UUID(64'd2559007593350444869 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_39 (.en(wire_7), .in(wire_24), .out(wire_43));
  TC_Switch # (.UUID(64'd4297414548625708919 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_40 (.en(wire_10), .in(wire_15), .out(wire_39));
  TC_Switch # (.UUID(64'd972928220399384192 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_41 (.en(wire_7), .in(wire_15), .out(wire_38));
  TC_Switch # (.UUID(64'd3044808667847191637 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_42 (.en(wire_10), .in(wire_35), .out(wire_58));
  TC_Switch # (.UUID(64'd2602597267482166209 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_43 (.en(wire_7), .in(wire_35), .out(wire_54));
  TC_Switch # (.UUID(64'd4266287403281139377 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_44 (.en(wire_10), .in(wire_52), .out(wire_46));
  TC_Switch # (.UUID(64'd1413005364500105444 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_45 (.en(wire_7), .in(wire_52), .out(wire_60));
  TC_Switch # (.UUID(64'd3142095426743800509 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_46 (.en(wire_10), .in(wire_26), .out(wire_27));
  TC_Switch # (.UUID(64'd793594983077177836 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_47 (.en(wire_7), .in(wire_26), .out(wire_31));
  TC_Register # (.UUID(64'd805183433895739842 ^ UUID), .BIT_WIDTH(64'd8)) Register8_48 (.clk(clk), .rst(rst), .load(wire_27), .save(wire_31), .in(wire_3), .out(wire_12_0));
  TC_Switch # (.UUID(64'd3523304946509383865 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_49 (.en(wire_10), .in(wire_28), .out(wire_36));
  TC_Switch # (.UUID(64'd3899091256447076266 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_50 (.en(wire_7), .in(wire_28), .out(wire_45));
  TC_Register # (.UUID(64'd197012223234376410 ^ UUID), .BIT_WIDTH(64'd8)) Register8_51 (.clk(clk), .rst(rst), .load(wire_36), .save(wire_45), .in(wire_3), .out(wire_12_2));
  TC_Switch # (.UUID(64'd1422811570386505738 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_52 (.en(wire_10), .in(wire_47), .out(wire_20));
  TC_Switch # (.UUID(64'd4182090768057833713 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_53 (.en(wire_7), .in(wire_47), .out(wire_29));
  TC_Register # (.UUID(64'd4311325631001493608 ^ UUID), .BIT_WIDTH(64'd8)) Register8_54 (.clk(clk), .rst(rst), .load(wire_20), .save(wire_29), .in(wire_3), .out(wire_12_5));
  TC_Switch # (.UUID(64'd3925860353481355705 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_55 (.en(wire_10), .in(wire_6), .out(wire_44));
  TC_Switch # (.UUID(64'd2354656880867171754 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_56 (.en(wire_7), .in(wire_6), .out(wire_0));
  TC_Register # (.UUID(64'd2497313757512643675 ^ UUID), .BIT_WIDTH(64'd8)) Register8_57 (.clk(clk), .rst(rst), .load(wire_44), .save(wire_0), .in(wire_3), .out(wire_12_7));
  _4bz_decoder # (.UUID(64'd4589577148535554959 ^ UUID)) _4bz_decoder_58 (.clk(clk), .rst(rst), .bit1(wire_55), .bit2(wire_61), .bit3(wire_11), .bit4(wire_34), .Disable(1'd0), .\8 (wire_24), .\9 (wire_15), .\10 (wire_52), .\11 (wire_35), .\12 (wire_28), .\13 (wire_26), .\14 (wire_47), .\15 (wire_6), .\0 (), .\1 (wire_32), .\2 (wire_30), .\3 (wire_1), .\4 (wire_17), .\5 (wire_40), .\6 (wire_4), .\7 (wire_13));
  TC_Constant # (.UUID(64'd4571590113858110367 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_59 (.out());
  TC_Constant # (.UUID(64'd3550419840356566641 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_60 (.out());

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  assign wire_2 = PUSH;
  wire [7:0] wire_3;
  assign wire_3 = VALUE;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  assign wire_5 = POP;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_12_0;
  wire [7:0] wire_12_1;
  wire [7:0] wire_12_2;
  wire [7:0] wire_12_3;
  wire [7:0] wire_12_4;
  wire [7:0] wire_12_5;
  wire [7:0] wire_12_6;
  wire [7:0] wire_12_7;
  wire [7:0] wire_12_8;
  wire [7:0] wire_12_9;
  wire [7:0] wire_12_10;
  wire [7:0] wire_12_11;
  wire [7:0] wire_12_12;
  wire [7:0] wire_12_13;
  wire [7:0] wire_12_14;
  assign wire_12 = wire_12_0|wire_12_1|wire_12_2|wire_12_3|wire_12_4|wire_12_5|wire_12_6|wire_12_7|wire_12_8|wire_12_9|wire_12_10|wire_12_11|wire_12_12|wire_12_13|wire_12_14;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_16_0;
  wire [7:0] wire_16_1;
  assign wire_16 = wire_16_0|wire_16_1;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_22_0;
  wire [0:0] wire_22_1;
  assign wire_22 = wire_22_0|wire_22_1;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [7:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;

endmodule
